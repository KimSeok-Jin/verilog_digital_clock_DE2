module OUTPUT(
    input TIMER_MODE,
    input ALARM_MODE,
    input SET_MODE,
    input SW_ACTIVE,
    input [3:0] TSEC0, TSEC1, TMIN0, TMIN1, THOUR0, THOUR1,
    input [3:0] ASEC0, ASEC1, AMIN0, AMIN1, AHOUR0, AHOUR1, ADAY0, ADAY1,
    input [3:0] SSEC0, SSEC1, SMIN0, SMIN1, SHOUR0, SHOUR1, SDAY0, SDAY1,
    input [3:0] SW_SEC0, SW_SEC1, SW_MIN0, SW_MIN1, SW_HOUR0, SW_HOUR1, SW_DAY0, SW_DAY1,
    input [3:0] SEC0, SEC1, MIN0, MIN1, HOUR0, HOUR1, DAY0, DAY1,
    output [3:0] OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7
);

    assign OUT0 = (TIMER_MODE) ? TSEC0 : (ALARM_MODE) ? ASEC0 : (SET_MODE) ? SSEC0 : (SW_ACTIVE) ? SW_SEC0 : SEC0;
    assign OUT1 = (TIMER_MODE) ? TSEC1 : (ALARM_MODE) ? ASEC1 : (SET_MODE) ? SSEC1 : (SW_ACTIVE) ? SW_SEC1 : SEC1;
    assign OUT2 = (TIMER_MODE) ? TMIN0 : (ALARM_MODE) ? AMIN0 : (SET_MODE) ? SMIN0 : (SW_ACTIVE) ? SW_MIN0 : MIN0;
    assign OUT3 = (TIMER_MODE) ? TMIN1 : (ALARM_MODE) ? AMIN1 : (SET_MODE) ? SMIN1 : (SW_ACTIVE) ? SW_MIN1 : MIN1;
    assign OUT4 = (TIMER_MODE) ? THOUR0 : (ALARM_MODE) ? AHOUR0 : (SET_MODE) ? SHOUR0 : (SW_ACTIVE) ? SW_HOUR0 : HOUR0;
    assign OUT5 = (TIMER_MODE) ? THOUR1 : (ALARM_MODE) ? AHOUR1 : (SET_MODE) ? SHOUR1 : (SW_ACTIVE) ? SW_HOUR1 : HOUR1;
    assign OUT6 = (TIMER_MODE) ? 4'b0000 : (ALARM_MODE) ? ADAY0 : (SET_MODE) ? SDAY0 : (SW_ACTIVE) ? SW_DAY0 : DAY0;
    assign OUT7 = (TIMER_MODE) ? 4'b0000 : (ALARM_MODE) ? ADAY1 : (SET_MODE) ? SDAY1 : (SW_ACTIVE) ? SW_DAY1 : DAY1;

endmodule 